library ieee;
use ieee.numeric_std.all;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

-- Author: Thomas Brown
-- Date: 11/13/19
-- Description: 2-bit counter that counts to 2.
entity count_to_two is
port (clk, reset, enable, enable_auto_reset : in std_logic;
      output : out std_logic_vector (1 downto 0));
end count_to_two;

architecture Behavioral of count_to_two is

signal temp_out : std_logic_vector (1 downto 0) := (others => '0');

begin

    process(clk, reset)
        begin
            if reset = '1' then
                temp_out <= (others => '0');
            elsif rising_edge(clk) then
                if enable = '1' then
                    if temp_out < 2 then
                        temp_out <= temp_out + 1;
                    elsif enable_auto_reset = '1' then
                        temp_out <= (others => '0');
                    end if;
                end if;
            end if;
        end process;

output <= temp_out;

end Behavioral;
